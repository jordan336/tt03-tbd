module jordan336_tbd (input [7:0] io_in,
                      output [7:0] io_out);
endmodule
